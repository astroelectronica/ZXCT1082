.title KiCad schematic
.include "C:/AE/ZXCT1082/_models/BZX84C4V7.spice.txt"
.include "C:/AE/ZXCT1082/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/ZXCT1082/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/ZXCT1082/_models/CGJ4C2C0G2A101J060AA_p.mod"
.include "C:/AE/ZXCT1082/_models/ZXCT1082.spice.txt"
R3 /PWR_IN /SP {RGT}
I1 /PWR_OUT 0 {ILOAD}
R2 /PWR_IN /PWR_OUT {RSENSE}
R1 /PWR_IN /PWR_OUT {RSENSE}
V1 /PWR_IN 0 {VSOURCE}
R4 /PWR_OUT /SN {RGT}
XU2 /SP /SN CGJ4C2C0G2A101J060AA_p
XU5 0 /OUT DI_BZX84C4V7
XU4 /OUT 0 C2012C0G2A102J060AA_p
R5 /COCM 0 {RG}
R6 /COCM /OUT {RLPF}
XU1 /COCM 0 /SP /SN VDD ZXCT1082
XU3 VDD 0 C2012X7R2A104K125AA_p
V2 VDD 0 {VSUPPLY}
.end
